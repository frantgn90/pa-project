
/*
 * This is the top level entity for the DECODE stage
 */

module decode_top();
	// Input signals

	// Output signals

	// Net type declaration

	// Port connections
endmodule